// An inferred RAM module of size 32x512
// Uses the ram512.mif file for its initial contents
module ram512(
	output reg [31:0] data_out,
	input wire [31:0] data_in, 
	input wire [8:0] address,
	input wire read, write
	
);

reg [31:0] i;

(*ram_file = "ram512.mif"*) reg [31:0] ram [0:511];

initial begin
	data_out = 32'b00000000000000000000000000000000;
	
//	// ORG $0
//	ram[0] <= 32'b00001_0011_0000_0000000000001010111; // ldi R3, $87
//	ram[1] <= 32'b00001_0011_0011_0000000000000000001; // ldi R3, 1(R3)
//	ram[2] <= 32'b00000_0010_0000_0000000000001000010; // ld R2, $66
//	ram[3] <= 32'b00001_0010_0010_1111111111111111111; // ldi R2, -1(R2)
//	ram[4] <= 32'b00011_0111_00000000000000000111101; // ldr R7, $61
//	ram[5] <= 32'b00100_0111_00000000000000000111100; // str $60, R7 ????
//	ram[6] <= 32'b00000_0001_0010_0000000000000000000; // ld R1, 0(R2)
//	ram[7] <= 32'b00001_0000_0000_0000000000000000001; // ldi R0, 1
//	ram[8] <= 32'b11011_000000000000000000000000000; // nop
//	ram[9] <= 32'b00101_0011_0010_0011_000000000000000; // add R3, R2, R3
//	ram[10] <= 32'b01101_0111_0111_0000000000000000010; // addi R7, R7, 2
//	ram[11] <= 32'b10010_0111_0111_0000000000000000000; // neg R7, R7
//	ram[12] <= 32'b10011_0111_0111_0000000000000000000; // not R7, R7
//	ram[13] <= 32'b01110_0111_0111_0000000000000001111; // andi R7, R7, $0F ??? Constant may be wrong
//	ram[14] <= 32'b01111_0111_0001_0000000000000000011; // ori R7, R1, 3
//	ram[15] <= 32'b01001_0010_0011_0000_000000000000000; // shr R2, R3, R0
//	ram[16] <= 32'b00010_0010_0000_0000000000000111000; // st $56, R2 ????
//	ram[17] <= 32'b01011_0001_0001_0000_000000000000000; // ror R1, R1, R0
//	ram[18] <= 32'b01100_0010_0010_0000_000000000000000; // rol R2, R2, R0
//	ram[19] <= 32'b01000_0010_0011_0000_000000000000000; // or R2, R3, R0
//	ram[20] <= 32'b00111_0001_0010_0001_000000000000000; // and R1, R2, R1
//	ram[21] <= 32'b00010_0011_0001_0000000000001001100; // st $4C(R1), R3 ???? (4C = 76)
//	ram[22] <= 32'b00110_0011_0010_0011_000000000000000; // sub R3, R2, R3
//	ram[23] <= 32'b01010_0001_0010_0000_000000000000000; // shl R1, R2, R0
//	ram[24] <= 32'b00001_0100_0000_0000000000000000101; // ldi R4, 5
//	ram[25] <= 32'b00001_0101_0000_0000000000000011111; // ldi R5, $1F (1F = 31)
//	ram[26] <= 32'b10000_0101_0100_0000000000000000000; // mul R5, R4
//	ram[27] <= 32'b11001_0111_00000000000000000000000; // mfhi R7
//	ram[28] <= 32'b11010_0110_00000000000000000000000; // mflo R6
//	ram[29] <= 32'b10001_0101_0100_0000000000000000000; // div R5, R4
//	ram[30] <= 32'b00001_1010_0100_0000000000000000000; // ldi R10, 0(R4)
//	ram[31] <= 32'b00001_1011_0101_0000000000000000000; // ldi R11, 0(R5)
//	ram[32] <= 32'b00001_1100_0110_0000000000000000000; // ldi R12, 0(R6)
//	ram[33] <= 32'b00001_1101_0111_0000000000000000000; // ldi R13, 0(R7)
//	ram[34] <= 32'b00001_1000_0000_0000000000000000100; // ldi R8, $4
//	ram[35] <= 32'b10110_1100_1110_0000000000000000100; // jal R12
//	ram[40] <= 32'b11101_1001_0000_0000000000000000000; // inc R9
//	ram[41] <= 32'b00001_0010_0000_0000000000000000011; // ldi R2, 3
//	ram[42] <= 32'b00001_0011_0000_0000000000000001010; // ldi R3, 10
//	ram[43] <= 32'b11100_000000000000000000000000000; // halt
//	
//	// ORG $9B
//	ram[155] <= 32'b11111_0100_0000_0000000000000000000; // ststk R4
//	ram[156] <= 32'b11111_1000_0000_0000000000000000000; // ststk R8
//	ram[157] <= 32'b00001_0100_0000_0000000000000001111; // ldi R4, $15
//	ram[158] <= 32'b00101_1001_1010_1100_000000000000000; // add R9, R10, R12
//	ram[159] <= 32'b00110_1000_1011_1101_000000000000000; // sub R8, R11, R13
//	ram[160] <= 32'b00110_1001_1001_1000_000000000000000; // sub R9, R9, R8
//	ram[161] <= 32'b11110_1000_0000_0000000000000000000; // ldstk R8
//	ram[162] <= 32'b11110_0100_0000_0000000000000000000; // ldstk R4
//	ram[163] <= 32'b10101_1110_00000000000000000000000; // jr R14
	
	ram[0] <= 32'b00001_0011_00000000000000000000110;
	ram[1] <= 32'b11111_0011_00000000000000000000000;
	ram[2] <= 32'b11101_0011_00000000000000000000000;
	ram[3] <= 32'b11110_0011_00000000000000000000000;
	ram[4] <= 32'b11100_000000000000000000000000000;

	// Values
	ram[66] <= 57;
	ram[56] <= 34;
	
end
	
always@(read, write) begin
	if(read == 1)
		data_out <= ram[address];
	else if(write == 1) begin
		ram[address] <= data_in;
		data_out <= 32'b00000000000000000000000000000000;
	end
	else
		data_out <= 32'b00000000000000000000000000000000;
end

endmodule
