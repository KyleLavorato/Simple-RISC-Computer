library verilog;
use verilog.vl_types.all;
entity Clock is
    port(
        clk             : out    vl_logic
    );
end Clock;
