library verilog;
use verilog.vl_types.all;
entity computerP3_tb is
end computerP3_tb;
